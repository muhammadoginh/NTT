`timescale 1ns / 1ps
`include "../rtl/Improved_Barrett_Reduction.v"
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/02/05 13:48:00
// Design Name: 
// Module Name: barrett2_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module barrett2_tb();

    // input
    reg clk;
    reg rstn;
    reg [95:0] X; // assumption X is a result of integer multiplication
    reg [47:0] q;
    reg [52:0] mu;
    
    // output
    wire [48:0] r;
    
    // instantiate unit under test
    barrett2 uut(
        .clk(clk),
        .rstn(rstn),
        .X(X),
        .q(q),
        .mu(mu),
        .r(r)
    );
    
    initial
    begin
        clk = 0;
        rstn = 1;
        q = 48'b111111111111111111111111111111111111110111110001;
        X = 96'b11101101110111001010010110110110111100010000001111101101110011000110010111110011000111011000;
        mu = 53'b01000000000000000000000000000000000000001000001111000;
        #1 rstn = 0;
        #9 X = 96'b1010001100000111001011011001000101000101100011100101001100000111111010110111010010001001110011;
            mu = 53'b1000000000000000000000000000000000000001000001111000;
        #10 X = 96'b10101001101011010000010111011000000000001001110111001010101100100000101100111000000110010010100;
            mu = 53'b1000000000000000000000000000000000000001000001111000;
        #10 X = 96'b1100110100000010011111000110000011011010111010101011110010100001011011010011010101010000100000;
            mu = 53'b1000000000000000000000000000000000000001000001111000;
        #10 X = 96'b1100110010011111101101010001001010110110011011010010110000000111101111100100101011110000110000;
            mu = 53'b1111111111111111111111111111111111111000001011100000;
            q = 48'b100000000000000000000000000000000000001111101001;
        #10 X = 96'b100001011000010011001010100011001001001100111101011110001010001111011101100111010001100011000;
            mu = 53'b1111111111111111111111111111111111111000001011100000;
        #10 X = 96'b1100100000111011101101111101110001111011000001010011001001000011101000100011110000000010000;
            mu = 53'b1111111111111111111111111111111111111000001011100000;
        #10 X = 96'b111011110011011111110100100001101100010001110010000010000101000000000010100110011110001110101;
            mu = 53'b1111111111111111111111111111111111111000001011100000;
    end
    
    always #1 clk = ~clk;
    
    initial $monitor("q=%b,X=%b,mu=%b,r=%b",q,X,mu,r);
    initial #80 $finish;
    
endmodule
